* Simple Circuit Example
V1 4 5 DC 10
V2 3 10 DC 5

R1 0 1 100
C1 1 2 100
R2 2 3 100
R3 0 4 200
R4 1 5 100
R5 2 6 100
R6 3 7 200
R7 4 5 100
C2 5 6 300
C3 6 7 100
R8 4 8 100
R9 5 9 200
R10 6 10 200
R11 7 11 300
C4 8 9 100
R12 9 10 200
R13 10 11 300

.tran 1ms 100ms
.control
run
plot V(1) V(2)
.endc
.end